// This is the unpowered netlist.
module tt_um_hsc_tdc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net15;
 wire net16;
 wire net2;
 wire net3;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire tdc_inst_capt_out_0 ;
 wire tdc_inst_capt_out_10 ;
 wire tdc_inst_capt_out_11 ;
 wire tdc_inst_capt_out_12 ;
 wire tdc_inst_capt_out_13 ;
 wire tdc_inst_capt_out_14 ;
 wire tdc_inst_capt_out_15 ;
 wire tdc_inst_capt_out_16 ;
 wire tdc_inst_capt_out_17 ;
 wire tdc_inst_capt_out_18 ;
 wire tdc_inst_capt_out_19 ;
 wire tdc_inst_capt_out_1 ;
 wire tdc_inst_capt_out_20 ;
 wire tdc_inst_capt_out_21 ;
 wire tdc_inst_capt_out_22 ;
 wire tdc_inst_capt_out_23 ;
 wire tdc_inst_capt_out_24 ;
 wire tdc_inst_capt_out_25 ;
 wire tdc_inst_capt_out_26 ;
 wire tdc_inst_capt_out_27 ;
 wire tdc_inst_capt_out_28 ;
 wire tdc_inst_capt_out_29 ;
 wire tdc_inst_capt_out_2 ;
 wire tdc_inst_capt_out_30 ;
 wire tdc_inst_capt_out_31 ;
 wire tdc_inst_capt_out_32 ;
 wire tdc_inst_capt_out_33 ;
 wire tdc_inst_capt_out_34 ;
 wire tdc_inst_capt_out_35 ;
 wire tdc_inst_capt_out_36 ;
 wire tdc_inst_capt_out_37 ;
 wire tdc_inst_capt_out_38 ;
 wire tdc_inst_capt_out_39 ;
 wire tdc_inst_capt_out_3 ;
 wire tdc_inst_capt_out_40 ;
 wire tdc_inst_capt_out_41 ;
 wire tdc_inst_capt_out_42 ;
 wire tdc_inst_capt_out_43 ;
 wire tdc_inst_capt_out_44 ;
 wire tdc_inst_capt_out_45 ;
 wire tdc_inst_capt_out_46 ;
 wire tdc_inst_capt_out_47 ;
 wire tdc_inst_capt_out_48 ;
 wire tdc_inst_capt_out_49 ;
 wire tdc_inst_capt_out_4 ;
 wire tdc_inst_capt_out_50 ;
 wire tdc_inst_capt_out_51 ;
 wire tdc_inst_capt_out_52 ;
 wire tdc_inst_capt_out_53 ;
 wire tdc_inst_capt_out_54 ;
 wire tdc_inst_capt_out_55 ;
 wire tdc_inst_capt_out_56 ;
 wire tdc_inst_capt_out_57 ;
 wire tdc_inst_capt_out_58 ;
 wire tdc_inst_capt_out_59 ;
 wire tdc_inst_capt_out_5 ;
 wire tdc_inst_capt_out_60 ;
 wire tdc_inst_capt_out_61 ;
 wire tdc_inst_capt_out_62 ;
 wire tdc_inst_capt_out_63 ;
 wire tdc_inst_capt_out_6 ;
 wire tdc_inst_capt_out_7 ;
 wire tdc_inst_capt_out_8 ;
 wire tdc_inst_capt_out_9 ;
 wire tdc_inst_capt_reg_r_1_0 ;
 wire tdc_inst_capt_reg_r_1_10 ;
 wire tdc_inst_capt_reg_r_1_11 ;
 wire tdc_inst_capt_reg_r_1_12 ;
 wire tdc_inst_capt_reg_r_1_13 ;
 wire tdc_inst_capt_reg_r_1_14 ;
 wire tdc_inst_capt_reg_r_1_15 ;
 wire tdc_inst_capt_reg_r_1_16 ;
 wire tdc_inst_capt_reg_r_1_17 ;
 wire tdc_inst_capt_reg_r_1_18 ;
 wire tdc_inst_capt_reg_r_1_19 ;
 wire tdc_inst_capt_reg_r_1_1 ;
 wire tdc_inst_capt_reg_r_1_20 ;
 wire tdc_inst_capt_reg_r_1_21 ;
 wire tdc_inst_capt_reg_r_1_22 ;
 wire tdc_inst_capt_reg_r_1_23 ;
 wire tdc_inst_capt_reg_r_1_24 ;
 wire tdc_inst_capt_reg_r_1_25 ;
 wire tdc_inst_capt_reg_r_1_26 ;
 wire tdc_inst_capt_reg_r_1_27 ;
 wire tdc_inst_capt_reg_r_1_28 ;
 wire tdc_inst_capt_reg_r_1_29 ;
 wire tdc_inst_capt_reg_r_1_2 ;
 wire tdc_inst_capt_reg_r_1_30 ;
 wire tdc_inst_capt_reg_r_1_31 ;
 wire tdc_inst_capt_reg_r_1_32 ;
 wire tdc_inst_capt_reg_r_1_33 ;
 wire tdc_inst_capt_reg_r_1_34 ;
 wire tdc_inst_capt_reg_r_1_35 ;
 wire tdc_inst_capt_reg_r_1_36 ;
 wire tdc_inst_capt_reg_r_1_37 ;
 wire tdc_inst_capt_reg_r_1_38 ;
 wire tdc_inst_capt_reg_r_1_39 ;
 wire tdc_inst_capt_reg_r_1_3 ;
 wire tdc_inst_capt_reg_r_1_40 ;
 wire tdc_inst_capt_reg_r_1_41 ;
 wire tdc_inst_capt_reg_r_1_42 ;
 wire tdc_inst_capt_reg_r_1_43 ;
 wire tdc_inst_capt_reg_r_1_44 ;
 wire tdc_inst_capt_reg_r_1_45 ;
 wire tdc_inst_capt_reg_r_1_46 ;
 wire tdc_inst_capt_reg_r_1_47 ;
 wire tdc_inst_capt_reg_r_1_48 ;
 wire tdc_inst_capt_reg_r_1_49 ;
 wire tdc_inst_capt_reg_r_1_4 ;
 wire tdc_inst_capt_reg_r_1_50 ;
 wire tdc_inst_capt_reg_r_1_51 ;
 wire tdc_inst_capt_reg_r_1_52 ;
 wire tdc_inst_capt_reg_r_1_53 ;
 wire tdc_inst_capt_reg_r_1_54 ;
 wire tdc_inst_capt_reg_r_1_55 ;
 wire tdc_inst_capt_reg_r_1_56 ;
 wire tdc_inst_capt_reg_r_1_57 ;
 wire tdc_inst_capt_reg_r_1_58 ;
 wire tdc_inst_capt_reg_r_1_59 ;
 wire tdc_inst_capt_reg_r_1_5 ;
 wire tdc_inst_capt_reg_r_1_60 ;
 wire tdc_inst_capt_reg_r_1_61 ;
 wire tdc_inst_capt_reg_r_1_62 ;
 wire tdc_inst_capt_reg_r_1_63 ;
 wire tdc_inst_capt_reg_r_1_6 ;
 wire tdc_inst_capt_reg_r_1_7 ;
 wire tdc_inst_capt_reg_r_1_8 ;
 wire tdc_inst_capt_reg_r_1_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_0 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_10 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_11 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_12 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_13 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_14 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_15 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_16 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_17 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_18 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_19 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_1 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_20 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_21 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_22 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_23 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_24 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_25 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_26 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_27 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_28 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_29 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_2 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_30 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_31 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_32 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_33 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_34 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_35 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_36 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_37 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_38 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_39 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_3 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_40 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_41 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_42 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_43 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_44 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_45 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_46 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_47 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_48 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_49 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_4 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_50 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_51 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_52 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_53 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_54 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_55 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_56 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_57 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_58 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_59 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_5 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_60 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_61 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_62 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_63 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_6 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_7 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_8 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_a_int_9 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_0 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_10 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_11 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_12 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_13 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_14 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_15 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_16 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_17 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_18 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_19 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_1 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_20 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_21 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_22 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_23 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_24 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_25 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_26 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_27 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_28 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_29 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_2 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_30 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_31 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_32 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_33 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_34 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_35 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_36 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_37 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_38 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_39 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_3 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_40 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_41 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_42 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_43 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_44 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_45 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_46 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_47 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_48 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_49 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_4 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_50 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_51 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_52 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_53 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_54 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_55 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_56 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_57 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_58 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_59 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_5 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_60 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_61 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_62 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_63 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_64 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_6 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_7 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_8 ;
 wire tdc_inst_dl_inst_dl_genblk_dl_ffout_w_9 ;
 wire tdc_inst_pc_inst_val_in ;
 wire tdc_inst_pc_inst_val_out ;
 wire tdc_inst_pg_pg_r_out ;
 wire tdc_inst_pg_val_r_out ;
 wire tdc_inst_pg_out ;
 wire tdc_inst_val_out_capt ;
 wire [1:0] clknet_0_ui_in;
 wire [0:0] clknet_1_0__leaf_ui_in;
 wire [0:0] clknet_1_1__leaf_ui_in;
 wire [1:0] clknet_4_0_0_ui_in;
 wire [1:0] clknet_4_10_0_ui_in;
 wire [1:0] clknet_4_11_0_ui_in;
 wire [1:0] clknet_4_12_0_ui_in;
 wire [1:0] clknet_4_13_0_ui_in;
 wire [1:0] clknet_4_14_0_ui_in;
 wire [1:0] clknet_4_15_0_ui_in;
 wire [1:0] clknet_4_1_0_ui_in;
 wire [1:0] clknet_4_2_0_ui_in;
 wire [1:0] clknet_4_3_0_ui_in;
 wire [1:0] clknet_4_4_0_ui_in;
 wire [1:0] clknet_4_5_0_ui_in;
 wire [1:0] clknet_4_6_0_ui_in;
 wire [1:0] clknet_4_7_0_ui_in;
 wire [1:0] clknet_4_8_0_ui_in;
 wire [1:0] clknet_4_9_0_ui_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(rst_n));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__mux2_1 _0470_ (.A0(net146),
    .A1(net5),
    .S(net3),
    .X(_0076_));
 sky130_fd_sc_hd__buf_1 _0471_ (.A(_0076_),
    .X(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_0 ));
 sky130_fd_sc_hd__inv_2 _0472_ (.A(net12),
    .Y(_0077_));
 sky130_fd_sc_hd__buf_2 _0473_ (.A(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0474_ (.A0(net4),
    .A1(net5),
    .S(net2),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_4 _0475_ (.A(net9),
    .X(_0080_));
 sky130_fd_sc_hd__or2_1 _0476_ (.A(_0080_),
    .B(net146),
    .X(_0081_));
 sky130_fd_sc_hd__buf_2 _0477_ (.A(rst_n),
    .X(_0082_));
 sky130_fd_sc_hd__buf_2 _0478_ (.A(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__o211a_1 _0479_ (.A1(_0078_),
    .A2(_0079_),
    .B1(_0081_),
    .C1(_0083_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_2 _0480_ (.A(_0080_),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _0481_ (.A(_0084_),
    .B(net33),
    .X(_0085_));
 sky130_fd_sc_hd__o211a_1 _0482_ (.A1(_0078_),
    .A2(net6),
    .B1(_0083_),
    .C1(_0085_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0483_ (.A0(net33),
    .A1(net6),
    .S(net3),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _0484_ (.A(_0080_),
    .B(tdc_inst_val_out_capt ),
    .X(_0087_));
 sky130_fd_sc_hd__o211a_1 _0485_ (.A1(_0078_),
    .A2(_0086_),
    .B1(_0087_),
    .C1(_0083_),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _0486_ (.A(_0084_),
    .B(tdc_inst_capt_reg_r_1_0 ),
    .X(_0088_));
 sky130_fd_sc_hd__o211a_1 _0487_ (.A1(_0078_),
    .A2(net83),
    .B1(_0083_),
    .C1(_0088_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _0488_ (.A(_0084_),
    .B(tdc_inst_capt_reg_r_1_1 ),
    .X(_0089_));
 sky130_fd_sc_hd__o211a_1 _0489_ (.A1(_0078_),
    .A2(net67),
    .B1(_0083_),
    .C1(_0089_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_2 _0490_ (.A(_0080_),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _0491_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_2 ),
    .X(_0091_));
 sky130_fd_sc_hd__o211a_1 _0492_ (.A1(_0078_),
    .A2(net70),
    .B1(_0083_),
    .C1(_0091_),
    .X(_0005_));
 sky130_fd_sc_hd__buf_2 _0493_ (.A(_0082_),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _0494_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_3 ),
    .X(_0093_));
 sky130_fd_sc_hd__o211a_1 _0495_ (.A1(_0078_),
    .A2(net77),
    .B1(_0092_),
    .C1(_0093_),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _0496_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_4 ),
    .X(_0094_));
 sky130_fd_sc_hd__o211a_1 _0497_ (.A1(_0078_),
    .A2(net45),
    .B1(_0092_),
    .C1(_0094_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _0498_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_5 ),
    .X(_0095_));
 sky130_fd_sc_hd__o211a_1 _0499_ (.A1(_0078_),
    .A2(net91),
    .B1(_0092_),
    .C1(_0095_),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _0500_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_6 ),
    .X(_0096_));
 sky130_fd_sc_hd__o211a_1 _0501_ (.A1(_0078_),
    .A2(net58),
    .B1(_0092_),
    .C1(_0096_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _0502_ (.A(_0077_),
    .X(_0097_));
 sky130_fd_sc_hd__or2_1 _0503_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_7 ),
    .X(_0098_));
 sky130_fd_sc_hd__o211a_1 _0504_ (.A1(_0097_),
    .A2(net65),
    .B1(_0092_),
    .C1(_0098_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _0505_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_8 ),
    .X(_0099_));
 sky130_fd_sc_hd__o211a_1 _0506_ (.A1(_0097_),
    .A2(net118),
    .B1(_0092_),
    .C1(_0099_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0507_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_9 ),
    .X(_0100_));
 sky130_fd_sc_hd__o211a_1 _0508_ (.A1(_0097_),
    .A2(net79),
    .B1(_0092_),
    .C1(_0100_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _0509_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_10 ),
    .X(_0101_));
 sky130_fd_sc_hd__o211a_1 _0510_ (.A1(_0097_),
    .A2(net110),
    .B1(_0092_),
    .C1(_0101_),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _0511_ (.A(_0090_),
    .B(tdc_inst_capt_reg_r_1_11 ),
    .X(_0102_));
 sky130_fd_sc_hd__o211a_1 _0512_ (.A1(_0097_),
    .A2(net39),
    .B1(_0092_),
    .C1(_0102_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_2 _0513_ (.A(net14),
    .X(_0103_));
 sky130_fd_sc_hd__or2_1 _0514_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_12 ),
    .X(_0104_));
 sky130_fd_sc_hd__o211a_1 _0515_ (.A1(_0097_),
    .A2(net60),
    .B1(_0092_),
    .C1(_0104_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_2 _0516_ (.A(_0082_),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _0517_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_13 ),
    .X(_0106_));
 sky130_fd_sc_hd__o211a_1 _0518_ (.A1(_0097_),
    .A2(net75),
    .B1(_0105_),
    .C1(_0106_),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _0519_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_14 ),
    .X(_0107_));
 sky130_fd_sc_hd__o211a_1 _0520_ (.A1(_0097_),
    .A2(net63),
    .B1(_0105_),
    .C1(_0107_),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _0521_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_15 ),
    .X(_0108_));
 sky130_fd_sc_hd__o211a_1 _0522_ (.A1(_0097_),
    .A2(net117),
    .B1(_0105_),
    .C1(_0108_),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _0523_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_16 ),
    .X(_0109_));
 sky130_fd_sc_hd__o211a_1 _0524_ (.A1(_0097_),
    .A2(net97),
    .B1(_0105_),
    .C1(_0109_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _0525_ (.A(_0077_),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _0526_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_17 ),
    .X(_0111_));
 sky130_fd_sc_hd__o211a_1 _0527_ (.A1(_0110_),
    .A2(net53),
    .B1(_0105_),
    .C1(_0111_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _0528_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_18 ),
    .X(_0112_));
 sky130_fd_sc_hd__o211a_1 _0529_ (.A1(_0110_),
    .A2(net106),
    .B1(_0105_),
    .C1(_0112_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _0530_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_19 ),
    .X(_0113_));
 sky130_fd_sc_hd__o211a_1 _0531_ (.A1(_0110_),
    .A2(net111),
    .B1(_0105_),
    .C1(_0113_),
    .X(_0022_));
 sky130_fd_sc_hd__or2_1 _0532_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_20 ),
    .X(_0114_));
 sky130_fd_sc_hd__o211a_1 _0533_ (.A1(_0110_),
    .A2(net47),
    .B1(_0105_),
    .C1(_0114_),
    .X(_0023_));
 sky130_fd_sc_hd__or2_1 _0534_ (.A(_0103_),
    .B(tdc_inst_capt_reg_r_1_21 ),
    .X(_0115_));
 sky130_fd_sc_hd__o211a_1 _0535_ (.A1(_0110_),
    .A2(net102),
    .B1(_0105_),
    .C1(_0115_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_2 _0536_ (.A(net13),
    .X(_0116_));
 sky130_fd_sc_hd__or2_1 _0537_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_22 ),
    .X(_0117_));
 sky130_fd_sc_hd__o211a_1 _0538_ (.A1(_0110_),
    .A2(net87),
    .B1(_0105_),
    .C1(_0117_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_2 _0539_ (.A(_0082_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_1 _0540_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_23 ),
    .X(_0119_));
 sky130_fd_sc_hd__o211a_1 _0541_ (.A1(_0110_),
    .A2(net56),
    .B1(_0118_),
    .C1(_0119_),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _0542_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_24 ),
    .X(_0120_));
 sky130_fd_sc_hd__o211a_1 _0543_ (.A1(_0110_),
    .A2(net72),
    .B1(_0118_),
    .C1(_0120_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _0544_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_25 ),
    .X(_0121_));
 sky130_fd_sc_hd__o211a_1 _0545_ (.A1(_0110_),
    .A2(net123),
    .B1(_0118_),
    .C1(_0121_),
    .X(_0028_));
 sky130_fd_sc_hd__or2_1 _0546_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_26 ),
    .X(_0122_));
 sky130_fd_sc_hd__o211a_1 _0547_ (.A1(_0110_),
    .A2(net61),
    .B1(_0118_),
    .C1(_0122_),
    .X(_0029_));
 sky130_fd_sc_hd__buf_2 _0548_ (.A(_0077_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _0549_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_27 ),
    .X(_0124_));
 sky130_fd_sc_hd__o211a_1 _0550_ (.A1(_0123_),
    .A2(net73),
    .B1(_0118_),
    .C1(_0124_),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _0551_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_28 ),
    .X(_0125_));
 sky130_fd_sc_hd__o211a_1 _0552_ (.A1(_0123_),
    .A2(net124),
    .B1(_0118_),
    .C1(_0125_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _0553_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_29 ),
    .X(_0126_));
 sky130_fd_sc_hd__o211a_1 _0554_ (.A1(_0123_),
    .A2(net43),
    .B1(_0118_),
    .C1(_0126_),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _0555_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_30 ),
    .X(_0127_));
 sky130_fd_sc_hd__o211a_1 _0556_ (.A1(_0123_),
    .A2(net51),
    .B1(_0118_),
    .C1(_0127_),
    .X(_0033_));
 sky130_fd_sc_hd__or2_1 _0557_ (.A(_0116_),
    .B(tdc_inst_capt_reg_r_1_31 ),
    .X(_0128_));
 sky130_fd_sc_hd__o211a_1 _0558_ (.A1(_0123_),
    .A2(net122),
    .B1(_0118_),
    .C1(_0128_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_2 _0559_ (.A(net12),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _0560_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_32 ),
    .X(_0130_));
 sky130_fd_sc_hd__o211a_1 _0561_ (.A1(_0123_),
    .A2(net69),
    .B1(_0118_),
    .C1(_0130_),
    .X(_0035_));
 sky130_fd_sc_hd__buf_2 _0562_ (.A(rst_n),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _0563_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_33 ),
    .X(_0132_));
 sky130_fd_sc_hd__o211a_1 _0564_ (.A1(_0123_),
    .A2(net132),
    .B1(_0131_),
    .C1(_0132_),
    .X(_0036_));
 sky130_fd_sc_hd__or2_1 _0565_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_34 ),
    .X(_0133_));
 sky130_fd_sc_hd__o211a_1 _0566_ (.A1(_0123_),
    .A2(net52),
    .B1(_0131_),
    .C1(_0133_),
    .X(_0037_));
 sky130_fd_sc_hd__or2_1 _0567_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_35 ),
    .X(_0134_));
 sky130_fd_sc_hd__o211a_1 _0568_ (.A1(_0123_),
    .A2(net137),
    .B1(_0131_),
    .C1(_0134_),
    .X(_0038_));
 sky130_fd_sc_hd__or2_1 _0569_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_36 ),
    .X(_0135_));
 sky130_fd_sc_hd__o211a_1 _0570_ (.A1(_0123_),
    .A2(net49),
    .B1(_0131_),
    .C1(_0135_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _0571_ (.A(_0077_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_1 _0572_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_37 ),
    .X(_0137_));
 sky130_fd_sc_hd__o211a_1 _0573_ (.A1(_0136_),
    .A2(net138),
    .B1(_0131_),
    .C1(_0137_),
    .X(_0040_));
 sky130_fd_sc_hd__or2_1 _0574_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_38 ),
    .X(_0138_));
 sky130_fd_sc_hd__o211a_1 _0575_ (.A1(_0136_),
    .A2(net37),
    .B1(_0131_),
    .C1(_0138_),
    .X(_0041_));
 sky130_fd_sc_hd__or2_1 _0576_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_39 ),
    .X(_0139_));
 sky130_fd_sc_hd__o211a_1 _0577_ (.A1(_0136_),
    .A2(net85),
    .B1(_0131_),
    .C1(_0139_),
    .X(_0042_));
 sky130_fd_sc_hd__or2_1 _0578_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_40 ),
    .X(_0140_));
 sky130_fd_sc_hd__o211a_1 _0579_ (.A1(_0136_),
    .A2(net36),
    .B1(_0131_),
    .C1(_0140_),
    .X(_0043_));
 sky130_fd_sc_hd__or2_1 _0580_ (.A(_0129_),
    .B(tdc_inst_capt_reg_r_1_41 ),
    .X(_0141_));
 sky130_fd_sc_hd__o211a_1 _0581_ (.A1(_0136_),
    .A2(net115),
    .B1(_0131_),
    .C1(_0141_),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_2 _0582_ (.A(net9),
    .X(_0142_));
 sky130_fd_sc_hd__or2_1 _0583_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_42 ),
    .X(_0143_));
 sky130_fd_sc_hd__o211a_1 _0584_ (.A1(_0136_),
    .A2(net35),
    .B1(_0131_),
    .C1(_0143_),
    .X(_0045_));
 sky130_fd_sc_hd__buf_2 _0585_ (.A(rst_n),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _0586_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_43 ),
    .X(_0145_));
 sky130_fd_sc_hd__o211a_1 _0587_ (.A1(_0136_),
    .A2(net130),
    .B1(_0144_),
    .C1(_0145_),
    .X(_0046_));
 sky130_fd_sc_hd__or2_1 _0588_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_44 ),
    .X(_0146_));
 sky130_fd_sc_hd__o211a_1 _0589_ (.A1(_0136_),
    .A2(net101),
    .B1(_0144_),
    .C1(_0146_),
    .X(_0047_));
 sky130_fd_sc_hd__or2_1 _0590_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_45 ),
    .X(_0147_));
 sky130_fd_sc_hd__o211a_1 _0591_ (.A1(_0136_),
    .A2(net55),
    .B1(_0144_),
    .C1(_0147_),
    .X(_0048_));
 sky130_fd_sc_hd__or2_1 _0592_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_46 ),
    .X(_0148_));
 sky130_fd_sc_hd__o211a_1 _0593_ (.A1(_0136_),
    .A2(net41),
    .B1(_0144_),
    .C1(_0148_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_2 _0594_ (.A(_0077_),
    .X(_0149_));
 sky130_fd_sc_hd__or2_1 _0595_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_47 ),
    .X(_0150_));
 sky130_fd_sc_hd__o211a_1 _0596_ (.A1(_0149_),
    .A2(net133),
    .B1(_0144_),
    .C1(_0150_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _0597_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_48 ),
    .X(_0151_));
 sky130_fd_sc_hd__o211a_1 _0598_ (.A1(_0149_),
    .A2(net144),
    .B1(_0144_),
    .C1(_0151_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _0599_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_49 ),
    .X(_0152_));
 sky130_fd_sc_hd__o211a_1 _0600_ (.A1(_0149_),
    .A2(net89),
    .B1(_0144_),
    .C1(_0152_),
    .X(_0052_));
 sky130_fd_sc_hd__or2_1 _0601_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_50 ),
    .X(_0153_));
 sky130_fd_sc_hd__o211a_1 _0602_ (.A1(_0149_),
    .A2(net140),
    .B1(_0144_),
    .C1(_0153_),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _0603_ (.A(_0142_),
    .B(tdc_inst_capt_reg_r_1_51 ),
    .X(_0154_));
 sky130_fd_sc_hd__o211a_1 _0604_ (.A1(_0149_),
    .A2(net108),
    .B1(_0144_),
    .C1(_0154_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_2 _0605_ (.A(net9),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _0606_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_52 ),
    .X(_0156_));
 sky130_fd_sc_hd__o211a_1 _0607_ (.A1(_0149_),
    .A2(net142),
    .B1(_0144_),
    .C1(_0156_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_2 _0608_ (.A(rst_n),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _0609_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_53 ),
    .X(_0158_));
 sky130_fd_sc_hd__o211a_1 _0610_ (.A1(_0149_),
    .A2(net120),
    .B1(_0157_),
    .C1(_0158_),
    .X(_0056_));
 sky130_fd_sc_hd__or2_1 _0611_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_54 ),
    .X(_0159_));
 sky130_fd_sc_hd__o211a_1 _0612_ (.A1(_0149_),
    .A2(net125),
    .B1(_0157_),
    .C1(_0159_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _0613_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_55 ),
    .X(_0160_));
 sky130_fd_sc_hd__o211a_1 _0614_ (.A1(_0149_),
    .A2(net81),
    .B1(_0157_),
    .C1(_0160_),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _0615_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_56 ),
    .X(_0161_));
 sky130_fd_sc_hd__o211a_1 _0616_ (.A1(_0149_),
    .A2(net127),
    .B1(_0157_),
    .C1(_0161_),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_4 _0617_ (.A(_0077_),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _0618_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_57 ),
    .X(_0163_));
 sky130_fd_sc_hd__o211a_1 _0619_ (.A1(_0162_),
    .A2(net93),
    .B1(_0157_),
    .C1(_0163_),
    .X(_0060_));
 sky130_fd_sc_hd__or2_1 _0620_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_58 ),
    .X(_0164_));
 sky130_fd_sc_hd__o211a_1 _0621_ (.A1(_0162_),
    .A2(net128),
    .B1(_0157_),
    .C1(_0164_),
    .X(_0061_));
 sky130_fd_sc_hd__or2_1 _0622_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_59 ),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _0623_ (.A1(_0162_),
    .A2(net99),
    .B1(_0157_),
    .C1(_0165_),
    .X(_0062_));
 sky130_fd_sc_hd__or2_1 _0624_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_60 ),
    .X(_0166_));
 sky130_fd_sc_hd__o211a_1 _0625_ (.A1(_0162_),
    .A2(net135),
    .B1(_0157_),
    .C1(_0166_),
    .X(_0063_));
 sky130_fd_sc_hd__or2_1 _0626_ (.A(_0155_),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0167_));
 sky130_fd_sc_hd__o211a_1 _0627_ (.A1(_0162_),
    .A2(net113),
    .B1(_0157_),
    .C1(_0167_),
    .X(_0064_));
 sky130_fd_sc_hd__or2_1 _0628_ (.A(_0080_),
    .B(tdc_inst_capt_reg_r_1_62 ),
    .X(_0168_));
 sky130_fd_sc_hd__o211a_1 _0629_ (.A1(_0162_),
    .A2(net104),
    .B1(_0157_),
    .C1(_0168_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_1 _0630_ (.A(_0080_),
    .B(net147),
    .X(_0169_));
 sky130_fd_sc_hd__o211a_1 _0631_ (.A1(_0162_),
    .A2(tdc_inst_capt_out_63 ),
    .B1(_0082_),
    .C1(_0169_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _0632_ (.A(tdc_inst_pc_inst_val_in ),
    .B(_0080_),
    .X(_0170_));
 sky130_fd_sc_hd__o211a_1 _0633_ (.A1(_0162_),
    .A2(net95),
    .B1(_0082_),
    .C1(_0170_),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _0634_ (.A(tdc_inst_capt_reg_r_1_60 ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(tdc_inst_capt_reg_r_1_43 ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _0636_ (.A(tdc_inst_capt_reg_r_1_58 ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(tdc_inst_capt_reg_r_1_54 ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(tdc_inst_capt_reg_r_1_50 ),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_1 _0639_ (.A(tdc_inst_capt_reg_r_1_26 ),
    .B(tdc_inst_capt_reg_r_1_22 ),
    .Y(_0176_));
 sky130_fd_sc_hd__or2_1 _0640_ (.A(tdc_inst_capt_reg_r_1_26 ),
    .B(tdc_inst_capt_reg_r_1_22 ),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _0641_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__xor2_1 _0642_ (.A(tdc_inst_capt_reg_r_1_32 ),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__inv_2 _0643_ (.A(tdc_inst_capt_reg_r_1_8 ),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _0644_ (.A(tdc_inst_capt_reg_r_1_63 ),
    .B(tdc_inst_capt_reg_r_1_14 ),
    .Y(_0181_));
 sky130_fd_sc_hd__or2_1 _0645_ (.A(tdc_inst_capt_reg_r_1_63 ),
    .B(tdc_inst_capt_reg_r_1_14 ),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _0646_ (.A(_0181_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__xor2_1 _0647_ (.A(tdc_inst_capt_reg_r_1_18 ),
    .B(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__xnor2_1 _0648_ (.A(_0180_),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__xor2_1 _0649_ (.A(_0179_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__xor2_2 _0650_ (.A(tdc_inst_capt_reg_r_1_33 ),
    .B(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_2 _0651_ (.A(tdc_inst_capt_reg_r_1_10 ),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _0652_ (.A(tdc_inst_capt_reg_r_1_41 ),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _0653_ (.A(tdc_inst_capt_reg_r_1_29 ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _0654_ (.A(tdc_inst_capt_reg_r_1_27 ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(tdc_inst_capt_reg_r_1_6 ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _0656_ (.A(tdc_inst_capt_reg_r_1_4 ),
    .Y(_0193_));
 sky130_fd_sc_hd__xor2_1 _0657_ (.A(tdc_inst_capt_reg_r_1_5 ),
    .B(tdc_inst_capt_reg_r_1_3 ),
    .X(_0194_));
 sky130_fd_sc_hd__xnor2_1 _0658_ (.A(tdc_inst_capt_reg_r_1_1 ),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__xnor2_1 _0659_ (.A(_0193_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__xnor2_1 _0660_ (.A(_0192_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__xnor2_1 _0661_ (.A(_0191_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__xnor2_1 _0662_ (.A(_0190_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__xnor2_1 _0663_ (.A(_0189_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__xor2_1 _0664_ (.A(_0188_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _0665_ (.A(tdc_inst_capt_reg_r_1_48 ),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__or2_1 _0666_ (.A(tdc_inst_capt_reg_r_1_48 ),
    .B(_0201_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_1 _0667_ (.A(_0202_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__xnor2_1 _0668_ (.A(_0175_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _0669_ (.A(tdc_inst_capt_reg_r_1_39 ),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _0670_ (.A(tdc_inst_capt_reg_r_1_37 ),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _0671_ (.A(tdc_inst_capt_reg_r_1_11 ),
    .B(tdc_inst_capt_reg_r_1_9 ),
    .Y(_0208_));
 sky130_fd_sc_hd__or2_1 _0672_ (.A(tdc_inst_capt_reg_r_1_11 ),
    .B(tdc_inst_capt_reg_r_1_9 ),
    .X(_0209_));
 sky130_fd_sc_hd__a21o_1 _0673_ (.A1(_0208_),
    .A2(_0209_),
    .B1(tdc_inst_capt_reg_r_1_7 ),
    .X(_0210_));
 sky130_fd_sc_hd__nand3_1 _0674_ (.A(tdc_inst_capt_reg_r_1_7 ),
    .B(_0208_),
    .C(_0209_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _0675_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(tdc_inst_capt_reg_r_1_2 ),
    .Y(_0213_));
 sky130_fd_sc_hd__xor2_1 _0677_ (.A(tdc_inst_capt_reg_r_1_21 ),
    .B(tdc_inst_capt_reg_r_1_17 ),
    .X(_0214_));
 sky130_fd_sc_hd__xnor2_1 _0678_ (.A(tdc_inst_capt_reg_r_1_13 ),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__xnor2_1 _0679_ (.A(_0213_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__or2_1 _0680_ (.A(_0212_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__nand2_1 _0681_ (.A(_0212_),
    .B(_0216_),
    .Y(_0218_));
 sky130_fd_sc_hd__and2_1 _0682_ (.A(_0217_),
    .B(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(tdc_inst_capt_reg_r_1_23 ),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(tdc_inst_capt_reg_r_1_0 ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(tdc_inst_capt_reg_r_1_47 ),
    .Y(_0222_));
 sky130_fd_sc_hd__xor2_1 _0686_ (.A(tdc_inst_capt_reg_r_1_31 ),
    .B(tdc_inst_capt_reg_r_1_28 ),
    .X(_0223_));
 sky130_fd_sc_hd__xnor2_1 _0687_ (.A(tdc_inst_capt_reg_r_1_25 ),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__xnor2_1 _0688_ (.A(_0222_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__xnor2_1 _0689_ (.A(_0221_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__xnor2_1 _0690_ (.A(_0220_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__xor2_1 _0691_ (.A(_0219_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__or2_1 _0692_ (.A(_0207_),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(_0207_),
    .B(_0228_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _0694_ (.A(_0229_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__xnor2_1 _0695_ (.A(_0206_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(tdc_inst_capt_reg_r_1_19 ),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _0697_ (.A(tdc_inst_capt_reg_r_1_38 ),
    .B(tdc_inst_capt_reg_r_1_36 ),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_1 _0698_ (.A(tdc_inst_capt_reg_r_1_38 ),
    .B(tdc_inst_capt_reg_r_1_36 ),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _0699_ (.A(_0234_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__xor2_2 _0700_ (.A(tdc_inst_capt_reg_r_1_34 ),
    .B(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(tdc_inst_capt_reg_r_1_16 ),
    .Y(_0238_));
 sky130_fd_sc_hd__xor2_2 _0702_ (.A(tdc_inst_capt_reg_r_1_44 ),
    .B(tdc_inst_capt_reg_r_1_42 ),
    .X(_0239_));
 sky130_fd_sc_hd__xnor2_2 _0703_ (.A(tdc_inst_capt_reg_r_1_40 ),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_2 _0704_ (.A(_0238_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__xor2_2 _0705_ (.A(_0237_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__xnor2_2 _0706_ (.A(tdc_inst_capt_reg_r_1_15 ),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_2 _0707_ (.A(_0233_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(tdc_inst_capt_reg_r_1_20 ),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(tdc_inst_capt_reg_r_1_24 ),
    .Y(_0246_));
 sky130_fd_sc_hd__xor2_1 _0710_ (.A(tdc_inst_capt_reg_r_1_51 ),
    .B(tdc_inst_capt_reg_r_1_49 ),
    .X(_0247_));
 sky130_fd_sc_hd__xnor2_1 _0711_ (.A(tdc_inst_capt_reg_r_1_46 ),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__xnor2_1 _0712_ (.A(_0246_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__xnor2_1 _0713_ (.A(_0245_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _0714_ (.A(tdc_inst_capt_reg_r_1_57 ),
    .B(tdc_inst_capt_reg_r_1_55 ),
    .Y(_0251_));
 sky130_fd_sc_hd__or2_1 _0715_ (.A(tdc_inst_capt_reg_r_1_57 ),
    .B(tdc_inst_capt_reg_r_1_55 ),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _0716_ (.A(_0251_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__xor2_1 _0717_ (.A(tdc_inst_capt_reg_r_1_53 ),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(tdc_inst_capt_reg_r_1_30 ),
    .Y(_0255_));
 sky130_fd_sc_hd__xor2_1 _0719_ (.A(tdc_inst_capt_reg_r_1_62 ),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0256_));
 sky130_fd_sc_hd__xnor2_1 _0720_ (.A(tdc_inst_capt_reg_r_1_59 ),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__xnor2_1 _0721_ (.A(_0255_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__xor2_1 _0722_ (.A(_0254_),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__xnor2_1 _0723_ (.A(tdc_inst_capt_reg_r_1_12 ),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__xor2_1 _0724_ (.A(_0250_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__xnor2_1 _0725_ (.A(tdc_inst_capt_reg_r_1_35 ),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__xor2_1 _0726_ (.A(_0244_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__xnor2_1 _0727_ (.A(tdc_inst_capt_reg_r_1_45 ),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__xor2_1 _0728_ (.A(_0232_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_1 _0729_ (.A(tdc_inst_capt_reg_r_1_52 ),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__xor2_1 _0730_ (.A(_0205_),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__xnor2_1 _0731_ (.A(tdc_inst_capt_reg_r_1_56 ),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__xnor2_1 _0732_ (.A(_0174_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__xnor2_1 _0733_ (.A(_0173_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__xnor2_1 _0734_ (.A(_0172_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__nor2_2 _0735_ (.A(_0171_),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__and2_1 _0736_ (.A(_0171_),
    .B(_0271_),
    .X(_0273_));
 sky130_fd_sc_hd__o21ai_1 _0737_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0084_),
    .Y(_0274_));
 sky130_fd_sc_hd__o211a_1 _0738_ (.A1(_0084_),
    .A2(uo_out[0]),
    .B1(_0082_),
    .C1(_0274_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _0739_ (.A(tdc_inst_capt_reg_r_1_33 ),
    .B(_0186_),
    .X(_0275_));
 sky130_fd_sc_hd__a21o_1 _0740_ (.A1(tdc_inst_capt_reg_r_1_10 ),
    .A2(_0187_),
    .B1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__o21ai_2 _0741_ (.A1(_0175_),
    .A2(_0204_),
    .B1(_0202_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_1 _0742_ (.A(_0189_),
    .B(_0199_),
    .X(_0278_));
 sky130_fd_sc_hd__o21a_1 _0743_ (.A1(_0188_),
    .A2(_0200_),
    .B1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__o21ai_1 _0744_ (.A1(_0206_),
    .A2(_0231_),
    .B1(_0229_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21bo_1 _0745_ (.A1(tdc_inst_capt_reg_r_1_32 ),
    .A2(_0177_),
    .B1_N(_0176_),
    .X(_0281_));
 sky130_fd_sc_hd__a21bo_1 _0746_ (.A1(tdc_inst_capt_reg_r_1_18 ),
    .A2(_0182_),
    .B1_N(_0181_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(_0180_),
    .B(_0184_),
    .X(_0283_));
 sky130_fd_sc_hd__o21a_1 _0748_ (.A1(_0179_),
    .A2(_0185_),
    .B1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__xnor2_1 _0749_ (.A(_0282_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__xor2_1 _0750_ (.A(_0281_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or2_1 _0751_ (.A(_0193_),
    .B(_0195_),
    .X(_0287_));
 sky130_fd_sc_hd__o21ai_2 _0752_ (.A1(_0192_),
    .A2(_0196_),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21a_1 _0753_ (.A1(_0213_),
    .A2(_0215_),
    .B1(_0217_),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(tdc_inst_capt_reg_r_1_5 ),
    .B(tdc_inst_capt_reg_r_1_3 ),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _0755_ (.A(tdc_inst_capt_reg_r_1_1 ),
    .B(_0194_),
    .Y(_0291_));
 sky130_fd_sc_hd__a22o_1 _0756_ (.A1(_0290_),
    .A2(_0291_),
    .B1(_0208_),
    .B2(_0211_),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__and4_1 _0758_ (.A(_0290_),
    .B(_0291_),
    .C(_0208_),
    .D(_0211_),
    .X(_0294_));
 sky130_fd_sc_hd__nor2_1 _0759_ (.A(_0293_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__xor2_1 _0760_ (.A(_0289_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__xor2_2 _0761_ (.A(_0288_),
    .B(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__or2_1 _0762_ (.A(_0191_),
    .B(_0197_),
    .X(_0298_));
 sky130_fd_sc_hd__o21a_1 _0763_ (.A1(_0190_),
    .A2(_0198_),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__xor2_1 _0764_ (.A(_0297_),
    .B(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__xnor2_1 _0765_ (.A(_0286_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_1 _0766_ (.A(_0280_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__xnor2_2 _0767_ (.A(_0279_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__or2_1 _0768_ (.A(_0220_),
    .B(_0226_),
    .X(_0304_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(_0227_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _0770_ (.A(_0219_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nand2_1 _0771_ (.A(tdc_inst_capt_reg_r_1_15 ),
    .B(_0242_),
    .Y(_0307_));
 sky130_fd_sc_hd__o21a_1 _0772_ (.A1(_0233_),
    .A2(_0243_),
    .B1(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__and2_1 _0773_ (.A(tdc_inst_capt_reg_r_1_21 ),
    .B(tdc_inst_capt_reg_r_1_17 ),
    .X(_0309_));
 sky130_fd_sc_hd__a21oi_1 _0774_ (.A1(tdc_inst_capt_reg_r_1_13 ),
    .A2(_0214_),
    .B1(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__a21boi_1 _0775_ (.A1(tdc_inst_capt_reg_r_1_34 ),
    .A2(_0235_),
    .B1_N(_0234_),
    .Y(_0311_));
 sky130_fd_sc_hd__and2_1 _0776_ (.A(tdc_inst_capt_reg_r_1_31 ),
    .B(tdc_inst_capt_reg_r_1_28 ),
    .X(_0312_));
 sky130_fd_sc_hd__a21oi_1 _0777_ (.A1(tdc_inst_capt_reg_r_1_25 ),
    .A2(_0223_),
    .B1(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(_0311_),
    .B(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _0779_ (.A(_0311_),
    .B(_0313_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_1 _0780_ (.A(_0314_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__or2_1 _0781_ (.A(_0222_),
    .B(_0224_),
    .X(_0317_));
 sky130_fd_sc_hd__o21a_1 _0782_ (.A1(_0221_),
    .A2(_0225_),
    .B1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__xnor2_1 _0783_ (.A(_0316_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__xnor2_1 _0784_ (.A(_0310_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__xnor2_1 _0785_ (.A(_0308_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21o_1 _0786_ (.A1(_0304_),
    .A2(_0306_),
    .B1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__nand3_1 _0787_ (.A(_0304_),
    .B(_0306_),
    .C(_0321_),
    .Y(_0323_));
 sky130_fd_sc_hd__and2_1 _0788_ (.A(_0322_),
    .B(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _0789_ (.A(_0238_),
    .B(_0240_),
    .X(_0325_));
 sky130_fd_sc_hd__o21a_1 _0790_ (.A1(_0237_),
    .A2(_0241_),
    .B1(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _0791_ (.A(_0246_),
    .B(_0248_),
    .X(_0327_));
 sky130_fd_sc_hd__o21a_1 _0792_ (.A1(_0245_),
    .A2(_0249_),
    .B1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__and2_1 _0793_ (.A(tdc_inst_capt_reg_r_1_44 ),
    .B(tdc_inst_capt_reg_r_1_42 ),
    .X(_0329_));
 sky130_fd_sc_hd__a21oi_1 _0794_ (.A1(tdc_inst_capt_reg_r_1_40 ),
    .A2(_0239_),
    .B1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xor2_1 _0795_ (.A(_0328_),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__xnor2_1 _0796_ (.A(_0326_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a21boi_1 _0797_ (.A1(tdc_inst_capt_reg_r_1_53 ),
    .A2(_0252_),
    .B1_N(_0251_),
    .Y(_0333_));
 sky130_fd_sc_hd__and2_1 _0798_ (.A(tdc_inst_capt_reg_r_1_51 ),
    .B(tdc_inst_capt_reg_r_1_49 ),
    .X(_0334_));
 sky130_fd_sc_hd__a21oi_1 _0799_ (.A1(tdc_inst_capt_reg_r_1_46 ),
    .A2(_0247_),
    .B1(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__or2_1 _0800_ (.A(_0333_),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0333_),
    .B(_0335_),
    .Y(_0337_));
 sky130_fd_sc_hd__and2_1 _0802_ (.A(_0336_),
    .B(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _0803_ (.A(tdc_inst_capt_reg_r_1_62 ),
    .B(tdc_inst_capt_reg_r_1_61 ),
    .X(_0339_));
 sky130_fd_sc_hd__a21o_1 _0804_ (.A1(tdc_inst_capt_reg_r_1_59 ),
    .A2(_0256_),
    .B1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _0805_ (.A(_0255_),
    .B(_0257_),
    .X(_0341_));
 sky130_fd_sc_hd__o21a_1 _0806_ (.A1(_0254_),
    .A2(_0258_),
    .B1(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__xnor2_1 _0807_ (.A(_0340_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__xnor2_1 _0808_ (.A(_0338_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _0809_ (.A(tdc_inst_capt_reg_r_1_12 ),
    .B(_0259_),
    .Y(_0345_));
 sky130_fd_sc_hd__o21a_1 _0810_ (.A1(_0250_),
    .A2(_0260_),
    .B1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__xor2_1 _0811_ (.A(_0344_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__xnor2_1 _0812_ (.A(_0332_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _0813_ (.A(tdc_inst_capt_reg_r_1_35 ),
    .B(_0261_),
    .Y(_0349_));
 sky130_fd_sc_hd__o21ai_1 _0814_ (.A1(_0244_),
    .A2(_0262_),
    .B1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__xnor2_1 _0815_ (.A(_0348_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__xnor2_1 _0816_ (.A(_0324_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(tdc_inst_capt_reg_r_1_45 ),
    .B(_0263_),
    .Y(_0353_));
 sky130_fd_sc_hd__o21ai_2 _0818_ (.A1(_0232_),
    .A2(_0264_),
    .B1(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__xnor2_2 _0819_ (.A(_0352_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__xnor2_2 _0820_ (.A(_0303_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(tdc_inst_capt_reg_r_1_52 ),
    .B(_0265_),
    .Y(_0357_));
 sky130_fd_sc_hd__o21a_1 _0822_ (.A1(_0205_),
    .A2(_0266_),
    .B1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__xor2_2 _0823_ (.A(_0356_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__xnor2_2 _0824_ (.A(_0277_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(tdc_inst_capt_reg_r_1_56 ),
    .B(_0267_),
    .Y(_0361_));
 sky130_fd_sc_hd__o21a_1 _0826_ (.A1(_0174_),
    .A2(_0268_),
    .B1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__xnor2_1 _0827_ (.A(_0360_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__xor2_1 _0828_ (.A(_0276_),
    .B(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(_0173_),
    .B(_0269_),
    .X(_0365_));
 sky130_fd_sc_hd__o21a_1 _0830_ (.A1(_0172_),
    .A2(_0270_),
    .B1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__xor2_1 _0831_ (.A(_0364_),
    .B(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__xor2_1 _0832_ (.A(_0272_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _0833_ (.A(_0080_),
    .B(uo_out[1]),
    .X(_0369_));
 sky130_fd_sc_hd__o211a_1 _0834_ (.A1(_0162_),
    .A2(_0368_),
    .B1(_0369_),
    .C1(_0083_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(_0360_),
    .B(_0362_),
    .X(_0370_));
 sky130_fd_sc_hd__or2b_1 _0836_ (.A(_0363_),
    .B_N(_0276_),
    .X(_0371_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(_0284_),
    .Y(_0372_));
 sky130_fd_sc_hd__and2_1 _0838_ (.A(_0281_),
    .B(_0285_),
    .X(_0373_));
 sky130_fd_sc_hd__a21o_1 _0839_ (.A1(_0282_),
    .A2(_0372_),
    .B1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__or2b_1 _0840_ (.A(_0301_),
    .B_N(_0280_),
    .X(_0375_));
 sky130_fd_sc_hd__or2b_1 _0841_ (.A(_0279_),
    .B_N(_0302_),
    .X(_0376_));
 sky130_fd_sc_hd__nand2_1 _0842_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _0843_ (.A(_0297_),
    .B(_0299_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21o_1 _0844_ (.A1(_0286_),
    .A2(_0300_),
    .B1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__o21ai_1 _0845_ (.A1(_0308_),
    .A2(_0320_),
    .B1(_0322_),
    .Y(_0380_));
 sky130_fd_sc_hd__o21ai_1 _0846_ (.A1(_0289_),
    .A2(_0294_),
    .B1(_0292_),
    .Y(_0381_));
 sky130_fd_sc_hd__or2b_1 _0847_ (.A(_0296_),
    .B_N(_0288_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(_0292_),
    .A1(_0381_),
    .S(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__xor2_1 _0849_ (.A(_0380_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__xor2_1 _0850_ (.A(_0379_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _0851_ (.A(_0316_),
    .B(_0318_),
    .X(_0386_));
 sky130_fd_sc_hd__o21ai_1 _0852_ (.A1(_0310_),
    .A2(_0319_),
    .B1(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__and2b_1 _0853_ (.A_N(_0326_),
    .B(_0331_),
    .X(_0388_));
 sky130_fd_sc_hd__o21ba_1 _0854_ (.A1(_0328_),
    .A2(_0330_),
    .B1_N(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__xnor2_1 _0855_ (.A(_0314_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__xnor2_1 _0856_ (.A(_0387_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(_0340_),
    .Y(_0392_));
 sky130_fd_sc_hd__or2_1 _0858_ (.A(_0392_),
    .B(_0342_),
    .X(_0393_));
 sky130_fd_sc_hd__a21boi_1 _0859_ (.A1(_0338_),
    .A2(_0343_),
    .B1_N(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__nor2_1 _0860_ (.A(_0336_),
    .B(_0393_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_1 _0861_ (.A1(_0336_),
    .A2(_0394_),
    .B1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_1 _0862_ (.A(_0344_),
    .B(_0346_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_1 _0863_ (.A1(_0332_),
    .A2(_0347_),
    .B1(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__xnor2_1 _0864_ (.A(_0396_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__xnor2_1 _0865_ (.A(_0391_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__or2b_1 _0866_ (.A(_0348_),
    .B_N(_0350_),
    .X(_0401_));
 sky130_fd_sc_hd__a21boi_1 _0867_ (.A1(_0324_),
    .A2(_0351_),
    .B1_N(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__xor2_1 _0868_ (.A(_0400_),
    .B(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__xnor2_1 _0869_ (.A(_0385_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__and2b_1 _0870_ (.A_N(_0352_),
    .B(_0354_),
    .X(_0405_));
 sky130_fd_sc_hd__a21oi_1 _0871_ (.A1(_0303_),
    .A2(_0355_),
    .B1(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__xnor2_1 _0872_ (.A(_0404_),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__xor2_1 _0873_ (.A(_0377_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_1 _0874_ (.A(_0356_),
    .B(_0358_),
    .Y(_0409_));
 sky130_fd_sc_hd__a21oi_1 _0875_ (.A1(_0277_),
    .A2(_0359_),
    .B1(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__xor2_1 _0876_ (.A(_0408_),
    .B(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__xnor2_1 _0877_ (.A(_0374_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__a21o_1 _0878_ (.A1(_0370_),
    .A2(_0371_),
    .B1(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__nand3_1 _0879_ (.A(_0370_),
    .B(_0371_),
    .C(_0412_),
    .Y(_0414_));
 sky130_fd_sc_hd__and2_1 _0880_ (.A(_0413_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_1 _0881_ (.A(_0364_),
    .B(_0366_),
    .Y(_0416_));
 sky130_fd_sc_hd__a21o_1 _0882_ (.A1(_0272_),
    .A2(_0367_),
    .B1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(_0415_),
    .B(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(_0415_),
    .B(_0417_),
    .Y(_0419_));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(_0418_),
    .B(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__or2_1 _0886_ (.A(_0080_),
    .B(uo_out[2]),
    .X(_0421_));
 sky130_fd_sc_hd__o211a_1 _0887_ (.A1(_0162_),
    .A2(_0420_),
    .B1(_0421_),
    .C1(_0083_),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _0888_ (.A(_0408_),
    .B(_0410_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _0889_ (.A(_0374_),
    .B(_0411_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _0890_ (.A(_0380_),
    .B(_0383_),
    .Y(_0424_));
 sky130_fd_sc_hd__a21bo_1 _0891_ (.A1(_0379_),
    .A2(_0384_),
    .B1_N(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__nor2_1 _0892_ (.A(_0292_),
    .B(_0382_),
    .Y(_0426_));
 sky130_fd_sc_hd__or2b_1 _0893_ (.A(_0390_),
    .B_N(_0387_),
    .X(_0427_));
 sky130_fd_sc_hd__o21a_1 _0894_ (.A1(_0314_),
    .A2(_0389_),
    .B1(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__xnor2_1 _0895_ (.A(_0426_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__and2_1 _0896_ (.A(_0391_),
    .B(_0399_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _0897_ (.A(_0395_),
    .B(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__and2b_1 _0898_ (.A_N(_0398_),
    .B(_0396_),
    .X(_0432_));
 sky130_fd_sc_hd__or3_1 _0899_ (.A(_0395_),
    .B(_0432_),
    .C(_0430_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _0900_ (.A(_0431_),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__xnor2_1 _0901_ (.A(_0429_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _0902_ (.A(_0400_),
    .B(_0402_),
    .Y(_0436_));
 sky130_fd_sc_hd__a21oi_1 _0903_ (.A1(_0385_),
    .A2(_0403_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__xnor2_1 _0904_ (.A(_0435_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__xor2_1 _0905_ (.A(_0425_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or2b_1 _0906_ (.A(_0407_),
    .B_N(_0377_),
    .X(_0440_));
 sky130_fd_sc_hd__o21a_1 _0907_ (.A1(_0404_),
    .A2(_0406_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__xnor2_1 _0908_ (.A(_0439_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_1 _0909_ (.A1(_0422_),
    .A2(_0423_),
    .B1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__and3_1 _0910_ (.A(_0422_),
    .B(_0423_),
    .C(_0442_),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_1 _0911_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a21oi_1 _0912_ (.A1(_0413_),
    .A2(_0419_),
    .B1(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__a31o_1 _0913_ (.A1(_0413_),
    .A2(_0419_),
    .A3(_0445_),
    .B1(_0077_),
    .X(_0447_));
 sky130_fd_sc_hd__o221a_1 _0914_ (.A1(_0084_),
    .A2(uo_out[3]),
    .B1(_0446_),
    .B2(_0447_),
    .C1(_0083_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _0915_ (.A(_0439_),
    .B(_0441_),
    .X(_0448_));
 sky130_fd_sc_hd__and2b_1 _0916_ (.A_N(_0438_),
    .B(_0425_),
    .X(_0449_));
 sky130_fd_sc_hd__o21bai_1 _0917_ (.A1(_0435_),
    .A2(_0437_),
    .B1_N(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21bo_1 _0918_ (.A1(_0429_),
    .A2(_0433_),
    .B1_N(_0431_),
    .X(_0451_));
 sky130_fd_sc_hd__or3_1 _0919_ (.A(_0292_),
    .B(_0382_),
    .C(_0428_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(_0431_),
    .A1(_0451_),
    .S(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__xnor2_1 _0921_ (.A(_0450_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(_0448_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__and2_1 _0923_ (.A(_0448_),
    .B(_0454_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(_0455_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__a21o_1 _0925_ (.A1(_0422_),
    .A2(_0423_),
    .B1(_0442_),
    .X(_0458_));
 sky130_fd_sc_hd__a21oi_1 _0926_ (.A1(_0413_),
    .A2(_0458_),
    .B1(_0444_),
    .Y(_0459_));
 sky130_fd_sc_hd__a31o_1 _0927_ (.A1(_0415_),
    .A2(_0417_),
    .A3(_0445_),
    .B1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__xnor2_1 _0928_ (.A(_0457_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_1 _0929_ (.A(_0084_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__o211a_1 _0930_ (.A1(_0084_),
    .A2(uo_out[4]),
    .B1(_0082_),
    .C1(_0462_),
    .X(_0072_));
 sky130_fd_sc_hd__and2b_1 _0931_ (.A_N(_0084_),
    .B(uo_out[5]),
    .X(_0463_));
 sky130_fd_sc_hd__o2bb2a_1 _0932_ (.A1_N(_0450_),
    .A2_N(_0453_),
    .B1(_0452_),
    .B2(_0431_),
    .X(_0464_));
 sky130_fd_sc_hd__a21oi_1 _0933_ (.A1(_0457_),
    .A2(_0460_),
    .B1(_0455_),
    .Y(_0465_));
 sky130_fd_sc_hd__o21ai_1 _0934_ (.A1(_0464_),
    .A2(_0465_),
    .B1(_0080_),
    .Y(_0466_));
 sky130_fd_sc_hd__a21oi_1 _0935_ (.A1(_0464_),
    .A2(_0465_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__o21a_1 _0936_ (.A1(_0463_),
    .A2(_0467_),
    .B1(_0083_),
    .X(_0073_));
 sky130_fd_sc_hd__o211a_1 _0937_ (.A1(_0084_),
    .A2(uo_out[6]),
    .B1(_0082_),
    .C1(_0466_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(tdc_inst_pc_inst_val_out ),
    .A1(tdc_inst_pc_inst_val_in ),
    .S(net15),
    .X(_0468_));
 sky130_fd_sc_hd__and2_1 _0939_ (.A(_0082_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _0940_ (.A(_0469_),
    .X(_0075_));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_1_1__leaf_ui_in[0]),
    .D(_0000_),
    .Q(tdc_inst_pg_pg_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_1_0__leaf_ui_in[0]),
    .D(_0001_),
    .Q(tdc_inst_pg_val_r_out ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(net34),
    .Q(tdc_inst_val_out_capt ));
 sky130_fd_sc_hd__dfxtp_1 _0944_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(net84),
    .Q(tdc_inst_capt_reg_r_1_0 ));
 sky130_fd_sc_hd__dfxtp_1 _0945_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net68),
    .Q(tdc_inst_capt_reg_r_1_1 ));
 sky130_fd_sc_hd__dfxtp_1 _0946_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net71),
    .Q(tdc_inst_capt_reg_r_1_2 ));
 sky130_fd_sc_hd__dfxtp_1 _0947_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net78),
    .Q(tdc_inst_capt_reg_r_1_3 ));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net46),
    .Q(tdc_inst_capt_reg_r_1_4 ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net92),
    .Q(tdc_inst_capt_reg_r_1_5 ));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net59),
    .Q(tdc_inst_capt_reg_r_1_6 ));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net66),
    .Q(tdc_inst_capt_reg_r_1_7 ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net119),
    .Q(tdc_inst_capt_reg_r_1_8 ));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(net80),
    .Q(tdc_inst_capt_reg_r_1_9 ));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0013_),
    .Q(tdc_inst_capt_reg_r_1_10 ));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net40),
    .Q(tdc_inst_capt_reg_r_1_11 ));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0015_),
    .Q(tdc_inst_capt_reg_r_1_12 ));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(net76),
    .Q(tdc_inst_capt_reg_r_1_13 ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(net64),
    .Q(tdc_inst_capt_reg_r_1_14 ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_4_13_0_ui_in[1]),
    .D(_0018_),
    .Q(tdc_inst_capt_reg_r_1_15 ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_4_11_0_ui_in[1]),
    .D(net98),
    .Q(tdc_inst_capt_reg_r_1_16 ));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net54),
    .Q(tdc_inst_capt_reg_r_1_17 ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net107),
    .Q(tdc_inst_capt_reg_r_1_18 ));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net112),
    .Q(tdc_inst_capt_reg_r_1_19 ));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net48),
    .Q(tdc_inst_capt_reg_r_1_20 ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net103),
    .Q(tdc_inst_capt_reg_r_1_21 ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net88),
    .Q(tdc_inst_capt_reg_r_1_22 ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net57),
    .Q(tdc_inst_capt_reg_r_1_23 ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(_0027_),
    .Q(tdc_inst_capt_reg_r_1_24 ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_4_8_0_ui_in[1]),
    .D(_0028_),
    .Q(tdc_inst_capt_reg_r_1_25 ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_4_9_0_ui_in[1]),
    .D(net62),
    .Q(tdc_inst_capt_reg_r_1_26 ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net74),
    .Q(tdc_inst_capt_reg_r_1_27 ));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_4_2_0_ui_in[1]),
    .D(_0031_),
    .Q(tdc_inst_capt_reg_r_1_28 ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(net44),
    .Q(tdc_inst_capt_reg_r_1_29 ));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0033_),
    .Q(tdc_inst_capt_reg_r_1_30 ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_4_2_0_ui_in[1]),
    .D(_0034_),
    .Q(tdc_inst_capt_reg_r_1_31 ));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0035_),
    .Q(tdc_inst_capt_reg_r_1_32 ));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0036_),
    .Q(tdc_inst_capt_reg_r_1_33 ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0037_),
    .Q(tdc_inst_capt_reg_r_1_34 ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(_0038_),
    .Q(tdc_inst_capt_reg_r_1_35 ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(net50),
    .Q(tdc_inst_capt_reg_r_1_36 ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net139),
    .Q(tdc_inst_capt_reg_r_1_37 ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(net38),
    .Q(tdc_inst_capt_reg_r_1_38 ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net86),
    .Q(tdc_inst_capt_reg_r_1_39 ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0043_),
    .Q(tdc_inst_capt_reg_r_1_40 ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_4_7_0_ui_in[1]),
    .D(net116),
    .Q(tdc_inst_capt_reg_r_1_41 ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_4_6_0_ui_in[1]),
    .D(_0045_),
    .Q(tdc_inst_capt_reg_r_1_42 ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net131),
    .Q(tdc_inst_capt_reg_r_1_43 ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0047_),
    .Q(tdc_inst_capt_reg_r_1_44 ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(_0048_),
    .Q(tdc_inst_capt_reg_r_1_45 ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net42),
    .Q(tdc_inst_capt_reg_r_1_46 ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net134),
    .Q(tdc_inst_capt_reg_r_1_47 ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net145),
    .Q(tdc_inst_capt_reg_r_1_48 ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net90),
    .Q(tdc_inst_capt_reg_r_1_49 ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net141),
    .Q(tdc_inst_capt_reg_r_1_50 ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net109),
    .Q(tdc_inst_capt_reg_r_1_51 ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net143),
    .Q(tdc_inst_capt_reg_r_1_52 ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_4_4_0_ui_in[1]),
    .D(net121),
    .Q(tdc_inst_capt_reg_r_1_53 ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net126),
    .Q(tdc_inst_capt_reg_r_1_54 ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net82),
    .Q(tdc_inst_capt_reg_r_1_55 ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(_0059_),
    .Q(tdc_inst_capt_reg_r_1_56 ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net94),
    .Q(tdc_inst_capt_reg_r_1_57 ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net129),
    .Q(tdc_inst_capt_reg_r_1_58 ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net100),
    .Q(tdc_inst_capt_reg_r_1_59 ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_5_0_ui_in[1]),
    .D(net136),
    .Q(tdc_inst_capt_reg_r_1_60 ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net114),
    .Q(tdc_inst_capt_reg_r_1_61 ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_1_0_ui_in[1]),
    .D(net105),
    .Q(tdc_inst_capt_reg_r_1_62 ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_4_12_0_ui_in[1]),
    .D(net148),
    .Q(tdc_inst_capt_reg_r_1_63 ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(net96),
    .Q(tdc_inst_pc_inst_val_in ));
 sky130_fd_sc_hd__dfxtp_2 _1009_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0068_),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_2 _1010_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0069_),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_2 _1011_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0070_),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_4 _1012_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0071_),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _1013_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0072_),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _1014_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0073_),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _1015_ (.CLK(clknet_4_15_0_ui_in[1]),
    .D(_0074_),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_4_14_0_ui_in[1]),
    .D(_0075_),
    .Q(tdc_inst_pc_inst_val_out ));
 sky130_fd_sc_hd__buf_2 _1033_ (.A(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_0 ),
    .X(tdc_inst_pg_out ));
 sky130_fd_sc_hd__buf_2 _1034_ (.A(tdc_inst_pc_inst_val_out ),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_ui_in_0  (.A(ui_in[0]),
    .X(clknet_0_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_ui_in_1  (.A(ui_in[1]),
    .X(clknet_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_ui_in_0  (.A(clknet_0_ui_in[0]),
    .X(clknet_1_0__leaf_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_ui_in_0  (.A(clknet_0_ui_in[0]),
    .X(clknet_1_1__leaf_ui_in[0]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_0_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_10_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_11_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_12_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_13_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_14_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_15_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_1_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_2_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_3_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_4_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_5_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_6_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_7_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_8_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_ui_in_1  (.A(clknet_0_ui_in[1]),
    .X(clknet_4_9_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net12),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net1),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net1),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net1),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net9),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(net12),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(tdc_inst_pg_val_r_out ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0049_),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(tdc_inst_capt_out_33 ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(tdc_inst_capt_out_47 ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0050_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(tdc_inst_capt_out_60 ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0063_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(tdc_inst_capt_out_35 ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(tdc_inst_capt_out_37 ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0040_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(tdc_inst_capt_out_50 ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0053_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(tdc_inst_capt_out_29 ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(tdc_inst_capt_out_52 ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0055_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(tdc_inst_capt_out_48 ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0051_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(tdc_inst_pg_pg_r_out ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(tdc_inst_capt_reg_r_1_63 ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0066_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0032_),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(tdc_inst_capt_out_4 ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0007_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(tdc_inst_capt_out_20 ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0023_),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(tdc_inst_capt_out_36 ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0039_),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(tdc_inst_capt_out_30 ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0002_),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(tdc_inst_capt_out_34 ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(tdc_inst_capt_out_17 ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0020_),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(tdc_inst_capt_out_45 ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(tdc_inst_capt_out_23 ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0026_),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(tdc_inst_capt_out_6 ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0009_),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(tdc_inst_capt_out_12 ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(tdc_inst_capt_out_26 ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(tdc_inst_capt_out_42 ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0029_),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(tdc_inst_capt_out_14 ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0017_),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(tdc_inst_capt_out_7 ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0010_),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(tdc_inst_capt_out_1 ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0004_),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(tdc_inst_capt_out_32 ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(tdc_inst_capt_out_2 ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0005_),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(tdc_inst_capt_out_40 ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(tdc_inst_capt_out_24 ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(tdc_inst_capt_out_27 ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0030_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(tdc_inst_capt_out_13 ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0016_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(tdc_inst_capt_out_3 ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0006_),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(tdc_inst_capt_out_9 ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0012_),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(tdc_inst_capt_out_55 ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(tdc_inst_capt_out_38 ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0058_),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(tdc_inst_capt_out_0 ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0003_),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(tdc_inst_capt_out_39 ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0042_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(tdc_inst_capt_out_22 ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0025_),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(tdc_inst_capt_out_49 ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0052_),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(tdc_inst_capt_out_5 ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0041_),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0008_),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(tdc_inst_capt_out_57 ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0060_),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(tdc_inst_val_out_capt ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0067_),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(tdc_inst_capt_out_16 ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0019_),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(tdc_inst_capt_out_59 ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0062_),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(tdc_inst_capt_out_44 ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(tdc_inst_capt_out_11 ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(tdc_inst_capt_out_21 ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0024_),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(tdc_inst_capt_out_62 ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0065_),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(tdc_inst_capt_out_18 ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0021_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(tdc_inst_capt_out_51 ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0054_),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(tdc_inst_capt_out_10 ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(tdc_inst_capt_out_19 ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0014_),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0022_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(tdc_inst_capt_out_61 ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0064_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(tdc_inst_capt_out_41 ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0044_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(tdc_inst_capt_out_15 ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(tdc_inst_capt_out_8 ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0011_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(tdc_inst_capt_out_53 ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0056_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(tdc_inst_capt_out_46 ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(tdc_inst_capt_out_31 ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(tdc_inst_capt_out_25 ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(tdc_inst_capt_out_28 ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(tdc_inst_capt_out_54 ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0057_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(tdc_inst_capt_out_56 ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(tdc_inst_capt_out_58 ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0061_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(tdc_inst_capt_out_43 ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0046_),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input1 (.A(ena),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_0_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_1 ),
    .DE(net16),
    .Q(tdc_inst_capt_out_0 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_10_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_11 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_10 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_11_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_12 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_11 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_12_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_13 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_12 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_13_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_14 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_13 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_14_DFE  (.CLK(clknet_4_11_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_15 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_14 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_15_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_16 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_15 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_16_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_17 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_16 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_17_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_18 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_17 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_18_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_19 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_18 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_19_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_20 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_19 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_1_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_2 ),
    .DE(net16),
    .Q(tdc_inst_capt_out_1 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_20_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_21 ),
    .DE(net14),
    .Q(tdc_inst_capt_out_20 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_21_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_22 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_21 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_22_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_23 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_22 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_23_DFE  (.CLK(clknet_4_9_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_24 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_23 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_24_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_25 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_24 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_25_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_26 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_25 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_26_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_27 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_26 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_27_DFE  (.CLK(clknet_4_8_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_28 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_27 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_28_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_29 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_28 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_29_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_30 ),
    .DE(net13),
    .Q(tdc_inst_capt_out_29 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_2_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_3 ),
    .DE(net16),
    .Q(tdc_inst_capt_out_2 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_30_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_31 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_30 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_31_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_32 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_31 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_32_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_33 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_32 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_33_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_34 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_33 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_34_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_35 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_34 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_35_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_36 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_35 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_36_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_37 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_36 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_37_DFE  (.CLK(clknet_4_2_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_38 ),
    .DE(net11),
    .Q(tdc_inst_capt_out_37 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_38_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_39 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_38 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_39_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_40 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_39 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_3_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_4 ),
    .DE(net16),
    .Q(tdc_inst_capt_out_3 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_40_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_41 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_40 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_41_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_42 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_41 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_42_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_43 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_42 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_43_DFE  (.CLK(clknet_4_6_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_44 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_43 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_44_DFE  (.CLK(clknet_4_6_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_45 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_44 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_45_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_46 ),
    .DE(net10),
    .Q(tdc_inst_capt_out_45 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_46_DFE  (.CLK(clknet_4_3_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_47 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_46 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_47_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_48 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_47 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_48_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_49 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_48 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_49_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_50 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_49 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_4_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_5 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_4 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_50_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_51 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_50 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_51_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_52 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_51 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_52_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_53 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_52 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_53_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_54 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_53 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_54_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_55 ),
    .DE(net8),
    .Q(tdc_inst_capt_out_54 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_55_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_56 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_55 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_56_DFE  (.CLK(clknet_4_1_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_57 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_56 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_57_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_58 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_57 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_58_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_59 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_58 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_59_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_60 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_59 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_5_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_6 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_5 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_60_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_61 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_60 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_61_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_62 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_61 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_62_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_63 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_62 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_63_DFE  (.CLK(clknet_4_0_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_64 ),
    .DE(net7),
    .Q(tdc_inst_capt_out_63 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_6_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_7 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_6 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_7_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_8 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_7 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_8_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_9 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_8 ));
 sky130_fd_sc_hd__edfxtp_1 tdc_inst_dl_capt_capt_genblk_9_DFE  (.CLK(clknet_4_10_0_ui_in[1]),
    .D(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_10 ),
    .DE(net15),
    .Q(tdc_inst_capt_out_9 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_0_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_0 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_0 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_1 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_10_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_10 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_10 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_11 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_11_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_11 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_11 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_12 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_12_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_12 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_12 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_13 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_13_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_13 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_13 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_14 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_14_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_14 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_14 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_15 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_15_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_15 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_15 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_16 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_16_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_16 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_16 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_17 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_17_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_17 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_17 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_18 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_18_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_18 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_18 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_19 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_19_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_19 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_19 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_20 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_1_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_1 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_1 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_2 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_20_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_20 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_20 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_21 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_21_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_21 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_21 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_22 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_22_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_22 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_22 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_23 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_23_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_23 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_23 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_24 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_24_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_24 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_24 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_25 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_25_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_25 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_25 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_26 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_26_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_26 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_26 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_27 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_27_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_27 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_27 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_28 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_28_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_28 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_28 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_29 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_29_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_29 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_29 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_30 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_2_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_2 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_2 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_3 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_30_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_30 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_30 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_31 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_31_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_31 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_31 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_32 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_32_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_32 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_32 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_33 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_33_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_33 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_33 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_34 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_34_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_34 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_34 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_35 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_35_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_35 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_35 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_36 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_36_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_36 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_36 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_37 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_37_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_37 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_37 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_38 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_38_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_38 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_38 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_39 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_39_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_39 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_39 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_40 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_3_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_3 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_3 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_4 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_40_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_40 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_40 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_41 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_41_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_41 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_41 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_42 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_42_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_42 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_42 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_43 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_43_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_43 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_43 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_44 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_44_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_44 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_44 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_45 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_45_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_45 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_45 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_46 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_46_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_46 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_46 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_47 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_47_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_47 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_47 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_48 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_48_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_48 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_48 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_49 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_49_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_49 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_49 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_50 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_4_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_4 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_4 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_5 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_50_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_50 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_50 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_51 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_51_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_51 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_51 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_52 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_52_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_52 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_52 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_53 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_53_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_53 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_53 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_54 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_54_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_54 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_54 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_55 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_55_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_55 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_55 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_56 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_56_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_56 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_56 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_57 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_57_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_57 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_57 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_58 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_58_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_58 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_58 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_59 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_59_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_59 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_59 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_60 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_5_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_5 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_5 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_6 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_60_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_60 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_60 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_61 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_61_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_61 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_61 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_62 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_62_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_62 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_62 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_63 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_63_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_63 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_63 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_64 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_6_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_6 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_6 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_7 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_7_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_7 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_7 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_8 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_8_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_8 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_8 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_9 ));
 sky130_fd_sc_hd__nand2_1 tdc_inst_dl_inst_dl_genblk_dl_dnand_genblk_9_DN  (.A(tdc_inst_dl_inst_dl_genblk_dl_a_int_9 ),
    .B(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_9 ),
    .Y(tdc_inst_dl_inst_dl_genblk_dl_ffout_w_10 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_0_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_0 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_10_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_10 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_11_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_11 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_12_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_12 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_13_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_13 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_14_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_14 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_15_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_15 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_16_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_16 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_17_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_17 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_18_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_18 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_19_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_19 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_1_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_1 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_20_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_20 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_21_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_21 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_22_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_22 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_23_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_23 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_24_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_24 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_25_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_25 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_26_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_26 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_27_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_27 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_28_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_28 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_29_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_29 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_2_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_2 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_30_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_30 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_31_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_31 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_32_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_32 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_33_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_33 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_34_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_34 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_35_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_35 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_36_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_36 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_37_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_37 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_38_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_38 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_39_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_39 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_3_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_3 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_40_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_40 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_41_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_41 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_42_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_42 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_43_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_43 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_44_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_44 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_45_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_45 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_46_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_46 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_47_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_47 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_48_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_48 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_49_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_49 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_4_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_4 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_50_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_50 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_51_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_51 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_52_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_52 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_53_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_53 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_54_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_54 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_55_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_55 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_56_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_56 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_57_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_57 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_58_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_58 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_59_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_59 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_5_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_5 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_60_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_60 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_61_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_61 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_62_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_62 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_63_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_63 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_6_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_6 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_7_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_7 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_8_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_8 ));
 sky130_fd_sc_hd__conb_1 tdc_inst_dl_inst_dl_genblk_dl_ones_const_ones_genblk_9_const_one  (.HI(tdc_inst_dl_inst_dl_genblk_dl_a_int_9 ));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_25 (.HI(net25));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_26 (.HI(net26));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_27 (.HI(net27));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_28 (.HI(net28));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_29 (.HI(net29));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_30 (.HI(net30));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_31 (.HI(net31));
 sky130_fd_sc_hd__conb_1 tt_um_hsc_tdc_32 (.HI(net32));
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

